module text_processing
