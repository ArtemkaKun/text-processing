module latin

// Maps accented letters to normal latin letters without diacrilics.
// Adapted from: http://web.archive.org/web/20120918093154/http://lehelk.com/2011/05/06/script-to-remove-diacritics/
const latin_character_to_diacritics_map = {
	// vfmt off
	'A':  ['A', 'Ⓐ', 'Ａ', 'À', 'Á', 'Â', 'Ầ', 'Ấ', 'Ẫ', 'Ẩ', 'Ã', 'Ā', 'Ă', 'Ằ', 'Ắ', 'Ẵ', 'Ẳ', 'Ȧ', 'Ǡ', 'Ä', 'Ǟ', 'Ả', 'Å', 'Ǻ', 'Ǎ', 'Ȁ', 'Ȃ', 'Ạ', 'Ậ', 'Ặ', 'Ḁ', 'Ą', 'Ⱥ', 'Ɐ']
	'AA': ['Ꜳ']
	'AE': ['Æ', 'Ǽ', 'Ǣ']
	'AO': ['Ꜵ']
	'AU': ['Ꜷ']
	'AV': ['Ꜹ', 'Ꜻ']
	'AY': ['Ꜽ']
	'B':  ['B', 'Ⓑ', 'Ｂ', 'Ḃ', 'Ḅ', 'Ḇ', 'Ƀ', 'Ƃ', 'Ɓ']
	'C':  ['C', 'Ⓒ', 'Ｃ', 'Ć', 'Ĉ', 'Ċ', 'Č', 'Ç', 'Ḉ', 'Ƈ', 'Ȼ', 'Ꜿ']
	'D':  ['D', 'Ⓓ', 'Ｄ', 'Ḋ', 'Ď', 'Ḍ', 'Ḑ', 'Ḓ', 'Ḏ', 'Đ', 'Ƌ', 'Ɗ', 'Ɖ', 'Ꝺ']
	'DZ': ['Ǳ', 'Ǆ']
	'Dz': ['ǲ', 'ǅ']
	'E':  ['E', 'Ⓔ', 'Ｅ', 'È', 'É', 'Ê', 'Ề', 'Ế', 'Ễ', 'Ể', 'Ẽ', 'Ē', 'Ḕ', 'Ḗ', 'Ĕ', 'Ė', 'Ë', 'Ẻ', 'Ě', 'Ȅ', 'Ȇ', 'Ẹ', 'Ệ', 'Ȩ', 'Ḝ', 'Ę', 'Ḙ', 'Ḛ', 'Ɛ', 'Ǝ']
	'F':  ['F', 'Ⓕ', 'Ｆ', 'Ḟ', 'Ƒ', 'Ꝼ']
	'G':  ['G', 'Ⓖ', 'Ｇ', 'Ǵ', 'Ĝ', 'Ḡ', 'Ğ', 'Ġ', 'Ǧ', 'Ģ', 'Ǥ', 'Ɠ', 'Ꞡ', 'Ᵹ', 'Ꝿ']
	'H':  ['H', 'Ⓗ', 'Ｈ', 'Ĥ', 'Ḣ', 'Ḧ', 'Ȟ', 'Ḥ', 'Ḩ', 'Ḫ', 'Ħ', 'Ⱨ', 'Ⱶ', 'Ɥ']
	'I':  ['I', 'Ⓘ', 'Ｉ', 'Ì', 'Í', 'Î', 'Ĩ', 'Ī', 'Ĭ', 'İ', 'Ï', 'Ḯ', 'Ỉ', 'Ǐ', 'Ȉ', 'Ȋ', 'Ị', 'Į', 'Ḭ', 'Ɨ']
	'J':  ['J', 'Ⓙ', 'Ｊ', 'Ĵ', 'Ɉ']
	'K':  ['K', 'Ⓚ', 'Ｋ', 'Ḱ', 'Ǩ', 'Ḳ', 'Ķ', 'Ḵ', 'Ƙ', 'Ⱪ', 'Ꝁ', 'Ꝃ', 'Ꝅ', 'Ꞣ']
	'L':  ['L', 'Ⓛ', 'Ｌ', 'Ŀ', 'Ĺ', 'Ľ', 'Ḷ', 'Ḹ', 'Ļ', 'Ḽ', 'Ḻ', 'Ł', 'Ƚ', 'Ɫ', 'Ⱡ', 'Ꝉ', 'Ꝇ', 'Ꞁ']
	'LJ': ['Ǉ']
	'Lj': ['ǈ']
	'M':  ['M', 'Ⓜ', 'Ｍ', 'Ḿ', 'Ṁ', 'Ṃ', 'Ɱ', 'Ɯ']
	'N':  ['N', 'Ⓝ', 'Ｎ', 'Ǹ', 'Ń', 'Ñ', 'Ṅ', 'Ň', 'Ṇ', 'Ņ', 'Ṋ', 'Ṉ', 'Ƞ', 'Ɲ', 'Ꞑ', 'Ꞥ']
	'NJ': ['Ǌ']
	'Nj': ['ǋ']
	'O':  ['O', 'Ⓞ', 'Ｏ', 'Ò', 'Ó', 'Ô', 'Ồ', 'Ố', 'Ỗ', 'Ổ', 'Õ', 'Ṍ', 'Ȭ', 'Ṏ', 'Ō', 'Ṑ', 'Ṓ', 'Ŏ', 'Ȯ', 'Ȱ', 'Ö', 'Ȫ', 'Ỏ', 'Ő', 'Ǒ', 'Ȍ', 'Ȏ', 'Ơ', 'Ờ', 'Ớ', 'Ỡ', 'Ở', 'Ợ', 'Ọ', 'Ộ', 'Ǭ', 'Ø', 'Ǿ', 'Ɔ', 'Ɵ', 'Ꝋ', 'Ꝍ']
	'OI': ['Ƣ']
	'OO': ['Ꝏ']
	'OU': ['Ȣ']
	'P':  ['P', 'Ⓟ', 'Ｐ', 'Ṕ', 'Ṗ', 'Ƥ', 'Ᵽ', 'Ꝑ', 'Ꝓ', 'Ꝕ']
	'Q':  ['Q', 'Ⓠ', 'Ｑ', 'Ꝗ', 'Ꝙ', 'Ɋ']
	'R':  ['R', 'Ⓡ', 'Ｒ', 'Ŕ', 'Ṙ', 'Ř', 'Ȑ', 'Ȓ', 'Ṛ', 'Ṝ', 'Ŗ', 'Ṟ', 'Ɍ', 'Ɽ', 'Ꝛ', 'Ꞧ', 'Ꞃ']
	'S':  ['S', 'Ⓢ', 'Ｓ', 'ẞ', 'Ś', 'Ṥ', 'Ŝ', 'Ṡ', 'Š', 'Ṧ', 'Ṣ', 'Ṩ', 'Ș', 'Ş', 'Ȿ', 'Ꞩ', 'Ꞅ']
	'T':  ['T', 'Ⓣ', 'Ｔ', 'Ṫ', 'Ť', 'Ṭ', 'Ț', 'Ţ', 'Ṱ', 'Ṯ', 'Ŧ', 'Ƭ', 'Ʈ', 'Ⱦ', 'Ꞇ']
	'TZ': ['Ꜩ']
	'U':  ['U', 'Ⓤ', 'Ｕ', 'Ù', 'Ú', 'Û', 'Ũ', 'Ṹ', 'Ū', 'Ṻ', 'Ŭ', 'Ü', 'Ǜ', 'Ǘ', 'Ǖ', 'Ǚ', 'Ủ', 'Ů', 'Ű', 'Ǔ', 'Ȕ', 'Ȗ', 'Ư', 'Ừ', 'Ứ', 'Ữ', 'Ử', 'Ự', 'Ụ', 'Ṳ', 'Ų', 'Ṷ', 'Ṵ', 'Ʉ']
	'V':  ['V', 'Ⓥ', 'Ｖ', 'Ṽ', 'Ṿ', 'Ʋ', 'Ꝟ', 'Ʌ']
	'VY': ['Ꝡ']
	'W':  ['W', 'Ⓦ', 'Ｗ', 'Ẁ', 'Ẃ', 'Ŵ', 'Ẇ', 'Ẅ', 'Ẉ', 'Ⱳ']
	'X':  ['X', 'Ⓧ', 'Ｘ', 'Ẋ', 'Ẍ']
	'Y':  ['Y', 'Ⓨ', 'Ｙ', 'Ỳ', 'Ý', 'Ŷ', 'Ỹ', 'Ȳ', 'Ẏ', 'Ÿ', 'Ỷ', 'Ỵ', 'Ƴ', 'Ɏ', 'Ỿ']
	'Z':  ['Z', 'Ⓩ', 'Ｚ', 'Ź', 'Ẑ', 'Ż', 'Ž', 'Ẓ', 'Ẕ', 'Ƶ', 'Ȥ', 'Ɀ', 'Ⱬ', 'Ꝣ']
	'a':  ['a', 'ⓐ', 'ａ', 'ẚ', 'à', 'á', 'â', 'ầ', 'ấ', 'ẫ', 'ẩ', 'ã', 'ā', 'ă', 'ằ', 'ắ', 'ẵ', 'ẳ', 'ȧ', 'ǡ', 'ä', 'ǟ', 'ả', 'å', 'ǻ', 'ǎ', 'ȁ', 'ȃ', 'ạ', 'ậ', 'ặ', 'ḁ', 'ą', 'ⱥ', 'ɐ']
	'aa': ['ꜳ']
	'ae': ['æ', 'ǽ', 'ǣ']
	'ao': ['ꜵ']
	'au': ['ꜷ']
	'av': ['ꜹ', 'ꜻ']
	'ay': ['ꜽ']
	'b':  ['b', 'ⓑ', 'ｂ', 'ḃ', 'ḅ', 'ḇ', 'ƀ', 'ƃ', 'ɓ']
	'c':  ['c', 'ⓒ', 'ｃ', 'ć', 'ĉ', 'ċ', 'č', 'ç', 'ḉ', 'ƈ', 'ȼ', 'ꜿ', 'ↄ']
	'd':  ['d', 'ⓓ', 'ｄ', 'ḋ', 'ď', 'ḍ', 'ḑ', 'ḓ', 'ḏ', 'đ', 'ƌ', 'ɖ', 'ɗ', 'ꝺ']
	'dz': ['ǳ', 'ǆ']
	'e':  ['e', 'ⓔ', 'ｅ', 'è', 'é', 'ê', 'ề', 'ế', 'ễ', 'ể', 'ẽ', 'ē', 'ḕ', 'ḗ', 'ĕ', 'ė', 'ë', 'ẻ', 'ě', 'ȅ', 'ȇ', 'ẹ', 'ệ', 'ȩ', 'ḝ', 'ę', 'ḙ', 'ḛ', 'ɇ', 'ɛ', 'ǝ']
	'f':  ['f', 'ⓕ', 'ｆ', 'ḟ', 'ƒ', 'ꝼ']
	'g':  ['g', 'ⓖ', 'ｇ', 'ǵ', 'ĝ', 'ḡ', 'ğ', 'ġ', 'ǧ', 'ģ', 'ǥ', 'ɠ', 'ꞡ', 'ᵹ', 'ꝿ']
	'h':  ['h', 'ⓗ', 'ｈ', 'ĥ', 'ḣ', 'ḧ', 'ȟ', 'ḥ', 'ḩ', 'ḫ', 'ẖ', 'ħ', 'ⱨ', 'ⱶ', 'ɥ']
	'hv': ['ƕ']
	'i':  ['i', 'ⓘ', 'ｉ', 'ì', 'í', 'î', 'ĩ', 'ī', 'ĭ', 'ï', 'ḯ', 'ỉ', 'ǐ', 'ȉ', 'ȋ', 'ị', 'į', 'ḭ', 'ɨ', 'ı']
	'j':  ['j', 'ⓙ', 'ｊ', 'ĵ', 'ǰ', 'ɉ']
	'k':  ['k', 'ⓚ', 'ｋ', 'ḱ', 'ǩ', 'ḳ', 'ķ', 'ḵ', 'ƙ', 'ⱪ', 'ꝁ', 'ꝃ', 'ꝅ', 'ꞣ']
	'l':  ['l', 'ⓛ', 'ｌ', 'ŀ', 'ĺ', 'ľ', 'ḷ', 'ḹ', 'ļ', 'ḽ', 'ḻ', 'ſ', 'ł', 'ƚ', 'ɫ', 'ⱡ', 'ꝉ', 'ꞁ', 'ꝇ']
	'lj': ['ǉ']
	'm':  ['m', 'ⓜ', 'ｍ', 'ḿ', 'ṁ', 'ṃ', 'ɱ', 'ɯ']
	'n':  ['n', 'ⓝ', 'ｎ', 'ǹ', 'ń', 'ñ', 'ṅ', 'ň', 'ṇ', 'ņ', 'ṋ', 'ṉ', 'ƞ', 'ɲ', 'ŉ', 'ꞑ', 'ꞥ']
	'nj': ['ǌ']
	'o':  ['o', 'ⓞ', 'ｏ', 'ò', 'ó', 'ô', 'ồ', 'ố', 'ỗ', 'ổ', 'õ', 'ṍ', 'ȭ', 'ṏ', 'ō', 'ṑ', 'ṓ', 'ŏ', 'ȯ', 'ȱ', 'ö', 'ȫ', 'ỏ', 'ő', 'ǒ', 'ȍ', 'ȏ', 'ơ', 'ờ', 'ớ', 'ỡ', 'ở', 'ợ', 'ọ', 'ộ', 'ǭ', 'ø', 'ǿ', 'ɔ', 'ꝋ', 'ꝍ', 'ɵ']
	'oi': ['ƣ']
	'ou': ['ȣ']
	'oo': ['ꝏ']
	'p':  ['p', 'ⓟ', 'ｐ', 'ṕ', 'ṗ', 'ƥ', 'ᵽ', 'ꝑ', 'ꝓ', 'ꝕ']
	'q':  ['q', 'ⓠ', 'ｑ', 'ɋ', 'ꝗ', 'ꝙ']
	'r':  ['r', 'ⓡ', 'ｒ', 'ŕ', 'ṙ', 'ř', 'ȑ', 'ȓ', 'ṛ', 'ṝ', 'ŗ', 'ṟ', 'ɍ', 'ɽ', 'ꝛ', 'ꞧ', 'ꞃ']
	's':  ['s', 'ⓢ', 'ｓ', 'ß', 'ś', 'ṥ', 'ŝ', 'ṡ', 'š', 'ṧ', 'ṣ', 'ṩ', 'ș', 'ş', 'ȿ', 'ꞩ', 'ꞅ', 'ẛ']
	't':  ['t', 'ⓣ', 'ｔ', 'ṫ', 'ẗ', 'ť', 'ṭ', 'ț', 'ţ', 'ṱ', 'ṯ', 'ŧ', 'ƭ', 'ʈ', 'ⱦ', 'ꞇ']
	'tz': ['ꜩ']
	'u':  ['u', 'ⓤ', 'ｕ', 'ù', 'ú', 'û', 'ũ', 'ṹ', 'ū', 'ṻ', 'ŭ', 'ü', 'ǜ', 'ǘ', 'ǖ', 'ǚ', 'ủ', 'ů', 'ű', 'ǔ', 'ȕ', 'ȗ', 'ư', 'ừ', 'ứ', 'ữ', 'ử', 'ự', 'ụ', 'ṳ', 'ų', 'ṷ', 'ṵ', 'ʉ']
	'v':  ['v', 'ⓥ', 'ｖ', 'ṽ', 'ṿ', 'ʋ', 'ꝟ', 'ʌ']
	'vy': ['ꝡ']
	'w':  ['w', 'ⓦ', 'ｗ', 'ẁ', 'ẃ', 'ŵ', 'ẇ', 'ẅ', 'ẘ', 'ẉ', 'ⱳ']
	'x':  ['x', 'ⓧ', 'ｘ', 'ẋ', 'ẍ']
	'y':  ['y', 'ⓨ', 'ｙ', 'ỳ', 'ý', 'ŷ', 'ỹ', 'ȳ', 'ẏ', 'ÿ', 'ỷ', 'ẙ', 'ỵ', 'ƴ', 'ɏ', 'ỿ']
	'z':  ['z', 'ⓩ', 'ｚ', 'ź', 'ẑ', 'ż', 'ž', 'ẓ', 'ẕ', 'ƶ', 'ȥ', 'ɀ', 'ⱬ', 'ꝣ']
	// vfmt on
}

// Returns a new string by exchanging the diacrylics of str by its latin counterparts,
// leaving untouched all other non Latin "characters".
pub fn normalize_latin_diacritics(str string) string {
	mut normalized_string := str.clone()

	for normalized_letter, characters_with_diacritics in latin.latin_character_to_diacritics_map {
		for character_with_diacritic in characters_with_diacritics {
			normalized_string = normalized_string.replace(character_with_diacritic, normalized_letter)
		}
	}

	return normalized_string
}
